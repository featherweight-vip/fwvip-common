
`ifndef INCLUDED_FWVIP_MACROS_SVH
`define INCLUDED_FWVIP_MACROS_SVH


`endif /* INCLUDED_FWVIP_MACROS_SVH */